library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.vcomponents.all;

-- Only XST supports RAM inference
-- Infers Single Port Block Ram

entity alu_mult_atpg_bram_hi is
    port(   clk : in  std_logic;
            we  : in  std_logic;
            en  : in  std_logic;
            ssr : in  std_logic;
            dop : out std_logic_vector(0 downto 0);
            a   : in  std_logic_vector(6 downto 0);
            di  : in  std_logic_vector(31 downto 0);
            do  : out std_logic_vector(31 downto 0));
end alu_mult_atpg_bram_hi;

-- 2K x 8 RAM Bank

architecture Structural of alu_mult_atpg_bram_hi is

begin

--    RAMB16_S9_inst : RAMB16_S9
--    generic map (
--        INIT => X"000",                 --  Value of output RAM registers at startup
--        SRVAL => X"000",                --  Ouput value upon SSR assertion
--        WRITE_MODE => "WRITE_FIRST",    --  WRITE_FIRST, READ_FIRST or NO_CHANGE
--
--        -- The following INIT_xx declarations specify the initial contents of the RAM
--
--        -- Address 0 to 511
--        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
--
--      -- Address 512 to 1023
--        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
--
--        -- Address 1024 to 1535
--        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
--
--        -- Address 1536 to 2047
--        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
--
--        -- The next set of INITP_xx are for the parity bits
--
--        -- Address 0 to 511
--        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--
--        -- Address 512 to 1023
--        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--
--        -- Address 1024 to 1535
--        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--
--        -- Address 1536 to 2047
--        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
--
--    port map (
--        DO      => do,              -- 8-bit Data Output
--        DOP     => dop,             -- Parity Output
--        ADDR    => a,               -- 11-bit Address Input
--        CLK     => clk,             -- Clock
--        DI      => di,              -- 8-bit Data Input
--        DIP     => di(7 downto 7),  -- Parity Input
--        EN      => en,              -- RAM Enable Input
--        SSR     => ssr,             -- Synchronous Set/Reset Input
--        WE      =>  we              -- Write Enable Input
--        );
--
--    -- End of RAMB16_S9_inst instantiation

end Structural;
