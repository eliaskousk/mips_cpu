library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity alu_mult_atpg_bram_lo is
    port(   clk         : in  std_logic;
            en          : in  std_logic;
            address     : in  std_logic_vector(6 downto 0);
            data_vector : out std_logic_vector(31 downto 0));
end alu_mult_atpg_bram_lo;

architecture Structural of alu_mult_atpg_bram_lo is

    type atpg_rom is array (0 to 127) of std_logic_vector(31 downto 0);

    constant vectors_lo: atpg_rom := (
        "00000000000000000000000000000000",
        "00000000001000100000000000000000",
        "10000100000000000000000001111111",
        "10100000110011100000000000000011",
        "10111101110101111100000001111100",
        "00000000000000000000110101000100",
        "00000111110001000000000000000110",
        "01111110000111110101110010011111",
        "01110100000000000001100000000000",
        "00000000000000000110000000010000",
        "11110010100111110011000011001000",
        "00001010000000000000110000000000",
        "00000000000000001101000000001110",
        "00000000000100111000100100001001",
        "00000000000000000100100000000111",
        "00000001100000000000000001111111",
        "00000000000000000000000000000101",
        "00110011011000000000001100000100",
        "00000110110100110100110010001001",
        "11010000000000000000000011000000",
        "00111010000000000000011000001000",
        "01101000000000000010000110000010",
        "00111000000011100000000000110010",
        "00000000000000000000000000011000",
        "11110000011000000000000000000000",
        "00100000000010000000001100000100",
        "00000000000000000000110000000100",
        "00000000000000000110000010100000",
        "01100100000000000000000000000100",
        "00000000000000000110000000000000",
        "11101000000000000000000000000000",
        "00000000000001110000100000010110",
        "10110100000100010000010000110010",
        "01010101110001110001011011100100",
        "11100011110100100000000000000000",
        "00000000110000000000000000000000",
        "00001001111000000000000000000110",
        "10000000000110000000001000010010",
        "11000010101001000000001000010010",
        "11011111000100010000011011001000",
        "01100110001000010000001100000100",
        "00000000000000000000010000001011",
        "10001100010001000001001011001000",
        "00100000000011101001000101001111",
        "11101000000000000000000000000000",
        "00000000000000000110111110111010",
        "10100000000010000110000000000010",
        "11010010011101001000000000000000",
        "10000101010000000000000110000010",
        "10100010000000111111001101000011",
        "00000011100000000000000000000101",
        "00100001100000000000000000000001",
        "01001001111001100001110000010010",
        "00000110010010010000000001111010",
        "11011000000000000000011000000000",
        "00000000000000011100111110000000",
        "10100000011000000001100000000100",
        "10010001111000000000000000000100",
        "00000000000000001000011000000001",
        "10100000000000000000000110000010",
        "10100000000000000000001100000100",
        "00000000000000000000110000010000",
        "00000000000000001100000000000000",
        "11101011001001000011000000001000",
        "00000000000000000001000000000001",
        "00010000000000001100101100111001",
        "11110000000000000000000000011000",
        "01110001001000000000000000000100",
        "00010000000000000000000001110010",
        "10000000000000110000000000000000",
        "11000000000000011000000000000000",
        "00000000000000000110000001001100",
        "00000101000000000011000000001000",
        "00001000000010000000000000000011",
        "11110110000000000000000011000000",
        "00100000001111000100000100110001",
        "00000100000000000000000001100000",
        "11111000000011000000000000001000",
        "00011000000000000000000001001100",
        "10000000010000110000000000010000",
        "00000000001100000000000000000000",
        "10000000000001001100000000010001",
        "00000000011000000000000000000100",
        "00000100010000001111100011110000",
        "00000000000000001000000000000001",
        "00000011110110010100110110000001",
        "00000000000000000000001000110010",
        "10000110000000000000010010110010",
        "00101000000011100000000000000000",
        "00001000111000000000000000000100",
        "00000000001000000010000000000110",
        "10001000100000000000000001000011",
        "11000000001000011000000000000001",
        "00110011000100001001001111001000",
        "11000110101100011100000001100100",
        "10001101011000110000000110000000",
        "00010000000110000000000000000000",
        "11100010000000001000000101100100",
        "00000000000000010000100010110010",
        "00000000001000000000000011001000",
        "01110000000100000000000000000011",
        "11100010110111010000110000000010",
        "10010001010100000000000000010101",
        "00001101000000000001000000001000",
        "00111010000000000010000110000010",
        "11010000000000000000000000000111",
        "00101000000000111110000111000011",
        "00000000000011100000000000000000",
        others => X"00000000");

begin

    process(clk, address)
    begin
        if(clk'event and clk = '1') then
            if en = '1' then
                data_vector <= vectors_lo(to_integer(unsigned(address)));
            else
                data_vector <= (others =>  '-');
            end if;
        end if;
    end process;

end Structural;
